library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--	In-Datapath-Out: Button endocoder and debounce => Pattern Encoder => 7seg Cathode Mux => 7seg endoder
	
--	Control: clock divider => Anode Sequencer & 7seg Cathode Mux == match anode and cathode to same digit

--	!!!!! USE SAME NAMES AS master_Lab1_Pt2.xdc for port IO !!!!!

entity Lab2_main is
    Port (	CLK100MHz: in std_logic;
			SW: in std_logic_vector(2 downto 0); -- use 3 switches as binary bits
			AN : out std_logic_vector(7 downto 0); --7 seg ANODES
			C : out std_logic_vector(7 downto 0) --7 seg Cathodes   order might be backward?
	);
end Lab2_main;

architecture Structural of Lab2_main is

	--Component Declarations:
	
	--ANDODE DECODER
	component AnnodeDecoder
	   Port (X: in std_logic_vector(2 downto 0); -- b bits "000" digCODE generated by clkDiv
		    AN_o: out std_logic_vector(7 downto 0)); --8 bits to select the annode to display on 
	end component;
		
	--PATTERN ENCODER
	component PatCoder
	Port (code : in STD_LOGIC_VECTOR (2 downto 0);	--input coded button push maybe better to just input the button?		
			pat_0 : out STD_LOGIC_VECTOR (4 downto 0);-- 4-1 bits 7seg character in hex, 0 bit for dot
			pat_1 : out STD_LOGIC_VECTOR (4 downto 0);
			pat_2 : out STD_LOGIC_VECTOR (4 downto 0);
			pat_3 : out STD_LOGIC_VECTOR (4 downto 0);
			pat_4 : out STD_LOGIC_VECTOR (4 downto 0);
			pat_5 : out STD_LOGIC_VECTOR (4 downto 0);
			pat_6 : out STD_LOGIC_VECTOR (4 downto 0);
			pat_7 : out STD_LOGIC_VECTOR (4 downto 0)
			);
	end component;
	
	--7SEG CATHODE MUX
	component Mux8to1_5bit
	Port (	I_0 : in std_logic_vector(4 downto 0); --4-1 bits are character, 0 bit is dot
			I_1 : in std_logic_vector(4 downto 0); -- 0 is dot on, 1 is dot off
			I_2 : in std_logic_vector(4 downto 0);
			I_3 : in std_logic_vector(4 downto 0);
			I_4 : in std_logic_vector(4 downto 0);
			I_5 : in std_logic_vector(4 downto 0);
			I_6 : in std_logic_vector(4 downto 0);
			I_7 : in std_logic_vector(4 downto 0);
			S : in  std_logic_vector(2 downto 0); --selection by clk div
			Z : out  std_logic_vector(4 downto 0) --out
			);  
	end component;
	
	--7SEG ENCODER
	component sevseg_dot
	Port ( int : in std_logic_vector (4 downto 1);--same input vector here
			dot : in std_logic;		--as here when using component. 4-1 bits are character in hex, 0 bit is dot
           seg : out std_logic_vector (7 downto 0));-- 7-1 bits are cathodes, 0 bit is dot. -- 0 is dot on, 1 is dot off	
	end component;

--signals for the interal wires connecting
signal clkdiv : std_logic_vector(10 downto 0); -- CLOCK 
signal digCode : std_logic_vector (2 downto 0); --signal from clock division for anode and cathode selection
--OBSOLETE signal btnCode : std_logic_vector (2 downto 0); --signal from buttons to pattern encoder to select the pattern
signal muxSegSig: std_logic_vector(4 downto 0); --signal from cathode mux to 7 seg encoder
signal pat_0,pat_1,pat_2,pat_3,pat_4,pat_5,pat_6,pat_7: std_logic_vector(4 downto 0);

begin
	clock_divider: process (CLK100MHz)		-- create system clock divder
	begin
		if (rising_edge(CLK100MHz)) then
			clkdiv <= clkdiv+1;
		end if;	    
	end process clock_divider;
	
	digit_select: process (clkdiv(10))
	begin
		if (rising_edge(clkdiv(10))) then
			case digCode is				--used to rotate 7 seg digits
		 		when "000" => digCode <= "001";
				when "001" => digCode <= "010";
				when "010" => digCode <= "011";
				when "011" => digCode <= "100";
				when "100" => digCode <= "101";
				when "101" => digCode <= "110";
				when "110" => digCode <= "111";
				when "111" => digCode <= "000";
			end case;
		end if;
	end process digit_select;
					
	PatternCoder: PatCoder port map(SW,pat_0,pat_1,pat_2,pat_3,pat_4,pat_5,pat_6,pat_7);
	--order of pat digits probably needs to flip, use anode selection. that's what enables the number anyway, or do it here
	
	--AnnodeDecoder
	ANdeCoder: AnnodeDecoder port map(digCode,AN); --I don't know if it'll let us output direct to AN hardware
		
	CathMux: Mux8to1_5bit port map(pat_0,pat_1,pat_2,pat_3,pat_4,pat_5,pat_6,pat_7,digcode,muxSegSig);--flip 7,6,5,4,3,2,1,0??
	CathCoder: sevseg_dot port map(muxSegSig,muxSegSig(0),C);

end Structural;
