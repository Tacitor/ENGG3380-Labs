-- VHDL code goes here